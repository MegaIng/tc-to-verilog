module TC_FullAdder (in0, in1, ci, out, co)
    input in0;
    input in1;
    input ci;
    output out;
    output co;
    
    assign out = in0 ^ in1 ^ ci;
    assign co = (in0 & in1) | ((in0 ^ in1) & ci);
endmodule

