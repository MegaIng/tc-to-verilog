module TC_Off(value);
    output value;
    
    assign value = 1'b0;
endmodule

