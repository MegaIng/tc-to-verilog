module TC_Or(a, b, out);
    input a;
    input b;
    output out;
    
    assign out = a | b;
endmodule

