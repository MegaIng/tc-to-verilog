module TC_Or3(in0, in1, in2, out);
    input in0;
    input in1;
    input in2;
    output out;
    
    assign out = in0 | in1 | in2;
endmodule

