module TC_On(value);
    output value;
    
    assign value = 1'b1;
endmodule

