module TC_Not(in, out);
    input in;
    output out;
       
    assign out = ~in;
endmodule

